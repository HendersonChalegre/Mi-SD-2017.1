`ifndef ALUOP
`define ALUOP

`define ALU_ADDU 4'd0 // 0000
`define ALU_SUBU 4'd1 // 0001
`define ALU_SLT  4'd2 // 0010
`define ALU_SLTU 4'd3 // 0011
`define ALU_AND  4'd4 // 0100
`define ALU_OR   4'd5 // 0101
`define ALU_XOR  4'd6 // 0110
`define ALU_LUI  4'd7 // 0111
`define ALU_SLL  4'd8 // 1000
`define ALU_SRL  4'd9 // 1001
`define ALU_SRA  4'd10 // 1010
`define ALU_NOR  4'd11 // 1011
`define ALU_XXX  4'd15 // 1100, 1101, 1110, 111	1

`endif //ALUOP

